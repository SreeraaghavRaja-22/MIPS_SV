module memory
#(parameter WIDTH = 32)
(
    input logic
)